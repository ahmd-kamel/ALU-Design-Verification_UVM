class alu_test extends uvm_test;

    `uvm_component_utils(alu_test)
    function new(string name = "alu_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction 
endclass